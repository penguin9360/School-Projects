// Complete the farmer module in this file
// Don't put any code in this file besides the farmer circuit

module farmer(e, f, x, g, b);

endmodule // farmer
