module farmer_test;

endmodule // farmer_test
